module ALU (
	input wire [31:0] input_1,
	input wire [31:0] input_2,
	input wire control,
	input wire reset);
endmodule