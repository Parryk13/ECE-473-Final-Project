// add


module add (
	input [31:0] NUMBER1, 
	input [31:0] NUMBER2, 
	output [31:0] SUM);

assign SUM = NUMBER1 + NUMBER2;

endmodule