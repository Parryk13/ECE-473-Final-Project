library verilog;
use verilog.vl_types.all;
entity registerarray_vlg_vec_tst is
end registerarray_vlg_vec_tst;
